`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:10:42 11/24/2016 
// Design Name:    chenyu
// Module Name:    DigitalClock 
// Project Name:   �����ܱ�
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DigitalClock(
    input rest,
    input start,
    input read
    );


endmodule
